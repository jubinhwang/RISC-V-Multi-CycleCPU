`timescale 1ns / 1ps

module ROM (
    input  logic [31:0] addr,
    output logic [31:0] data
);
    logic [31:0] rom[0:2**8-1];

    initial begin
        $readmemh("code.mem",rom);
        // **RISC-V RV32I R-Type 검증** 
        //초기값 x[i] = i
        /*
        // 1. ADD: x10 = x1 + x2
        // 예상 결과: x10 = 1 + 2 = 3
        rom[0] = 32'b0000000_00010_00001_000_01010_0110011;

        // 2. SUB: x11 = x4 - x3
        // 예상 결과: x11 = 4 - 3 = 1
        rom[1] = 32'b0100000_00011_00100_000_01011_0110011;

        // 3. XOR: x12 = x5 ^ x6
        // 예상 결과: x12 = 5 ^ 6 = 3
        rom[2] = 32'b0000000_00110_00101_100_01100_0110011;

        // 4. OR: x13 = x7 | x8
        // 예상 결과: x13 = 7 | 8 = 15
        rom[3] = 32'b0000000_01000_00111_110_01101_0110011;

        // 5. AND: x14 = x9 & x10 (x10은 rom[0]의 결과인 3)
        // 예상 결과: x14 = 9 & 3 = 1
        rom[4] = 32'b0000000_01010_01001_111_01110_0110011;

        // 6. SLL: x15 = x11 << x2 (x11은 rom[1]의 결과인 1)
        // 예상 결과: x15 = 1 << 2 = 4
        rom[5] = 32'b0000000_00010_01011_001_01111_0110011;

        // 7. SRL: x16 = x13 >> x3 (x13은 rom[3]의 결과인 15)
        // 예상 결과: x16 = 15 >> 3 = 1
        rom[6] = 32'b0000000_00011_01101_101_10000_0110011;
        
        // 8. SRA: x17 = x20 >> x4 
        // 예상 결과: x17 = 20 >> 4 = 1
        rom[7] = 32'b0100000_00100_10100_101_10001_0110011;

        // 9. SLT: x18 = x21 < x22 
        // 예상 결과: 21 < 22는 참이므로 x18 = 1
        rom[8] = 32'b0000000_10110_10101_010_10010_0110011;

        // 10. SLTU: x19 = x23 < x22 
        // 예상 결과: 23 < 22는 거짓이므로 x19 = 0
        rom[9] = 32'b0000000_10110_10111_011_10011_0110011;

        // 11. 테스트 종료 후 현재 위치로 무한 점프
        rom[10] = 32'h0000006F; // jal x0, 0
        */
        /*
        // **RISC-V RV32I I-Type 검증** 
        //초기값 x[i] = i
        // //rom[x]=32'b   imm      _ rs1 _ f3_ rd  _ opcode; // I-Type
        // --- I-Type : 산술 연산 (Arithmetic) ---
        // 1. ADDI: x8 = x1 + 10
        // 예상 결과: x8 = 1 + 10 = 11
        rom[0] = 32'b000000001010_00001_000_01000_0010011;

        // 2. SLTI: x9 = (x2 < 5) ? 1 : 0 (Signed)
        // 예상 결과: 2 < 5 는 참이므로 x9 = 1
        rom[1] = 32'b000000000101_00010_010_01001_0010011;

        // 3. SLTIU: x10 = (x3 < 2) ? 1 : 0 (Unsigned)
        // 예상 결과: 3 < 2 는 거짓이므로 x10 = 0
        rom[2] = 32'b000000000010_00011_011_01010_0010011;

        // --- I-Type : 논리 연산 (Logical) ---
        // 4. XORI: x11 = x3 ^ 15
        // 예상 결과: x11 = 3 (0b0011) ^ 15 (0b1111) = 12 (0b1100)
        rom[3] = 32'b000000001111_00011_100_01011_0010011;

        // 5. ORI: x12 = x5 | 8
        // 예상 결과: x12 = 5 (0b0101) | 8 (0b1000) = 13 (0b1101)
        rom[4] = 32'b000000001000_00101_110_01100_0010011;

        // 6. ANDI: x13 = x6 & 7
        // 예상 결과: x13 = 6 (0b0110) & 7 (0b0111) = 6 (0b0110)
        rom[5] = 32'b000000000111_00110_111_01101_0010011;

        // --- I-Type : 시프트 연산 (Shift) ---
        // 7. SLLI: x14 = x7 << 3 (shamt = 3)
        // 예상 결과: x14 = 7 << 3 = 56
        rom[6] = 32'b0000000_00011_00111_001_01110_0010011;

        // 8. SRLI: x15 = x9 >> 2 (shamt = 2)
        // 예상 결과: x15 = 9 >> 2 = 2
        rom[7] = 32'b0000000_00010_01001_101_01111_0010011;

        // 9. SRAI: x16 = x1 + (-2)  -> 먼저 x16 = -1 (0xFFFFFFFF) 만들기
        //          x17 = x16 >> 2 (shamt = 2)
        rom[8] = 32'b111111111110_00001_000_10000_0010011; // addi x16, x1, -2 (x16 = 1 + (-2) = -1)
        // 예상 결과 (SRAI): x17 = -1 >> 2 = -1 (0xFFFFFFFF) (부호 비트 유지)
        rom[9] = 32'b0100000_00010_10000_101_10001_0010011; // srai x17, x16, 2

        // rom[0] = 32'b000000000001_00001_000_01001_0010011;// addi x9, x1, 1;
        // rom[1] = 32'b000000000100_00010_111_01010_0010011;// andi x10, x2, 4;
        // rom[2] = 32'b000000000011_00001_001_01011_0010011;// slli x11, x1, 3;
        // rom[3] = 32'b000000001001_00001_001_01100_0010011;// slli x12, x1, 9;
        // rom[4] = 32'b000000011110_00001_001_01101_0010011;// slli x13, x1, 30;
        */

        /*
        // B-Type: imm[12,10:5] _ rs2 _ rs1 _ f3 _ imm[4:1,11] _ opcode
        // B-Type: imm[12,10:5] _ rs2 _ rs1 _ f3 _ imm[4:1,11] _ opcode
        // 모든 점프 offset은 8 (명령어 2개 분량)로 통일합니다.
        
        // --- 1. BNE (Taken) ---
        // [PC=0] rom[0]: bne x1, x2, 8 (x1 != x2 -> 참)
        // 분기 성공 위치: PC+8 = 8 (rom[2])
        rom[0] = 32'b0000000_00010_00001_001_01000_1100011;

        // --- 2. BLT (Taken) ---
        // [PC=8] rom[2]: blt x1, x2, 8 (x1 < x2 -> 참)
        // 분기 성공 위치: PC+8 = 16 (rom[4])
        rom[2] = 32'b0000000_00010_00001_100_01000_1100011;

        // --- 3. BLTU (Taken) ---
        // [PC=16] rom[4]: bltu x1, x2, 8 (x1 < x2 -> 참)
        // 분기 성공 위치: PC+8 = 24 (rom[6])
        rom[4] = 32'b0000000_00010_00001_110_01000_1100011;

        // --- 4. BGE (Taken) ---
        // [PC=24] rom[6]: bge x2, x1, 8 (x2 >= x1 -> 참)
        // 분기 성공 위치: PC+8 = 32 (rom[8])
        rom[6] = 32'b0000000_00001_00010_101_01000_1100011;

        // --- 5. BGEU (Taken) ---
        // [PC=32] rom[8]: bgeu x2, x1, 8 (x2 >= x1 -> 참)
        // 분기 성공 위치: PC+8 = 40 (rom[10])
        rom[8] = 32'b0000000_00001_00010_111_01000_1100011;

        // --- 6. BEQ (Taken) ---
        // [PC=40] rom[10]: beq x0, x0, 8 (x0 == x0 -> 참)
        // 분기 성공 위치: PC+8 = 48 (rom[12])
        rom[10] = 32'b0000000_00000_00000_000_01000_1100011;

        // --- 테스트 종료 ---
        // [PC=48] rom[12]: 무한 루프
        rom[12] = 32'h0000006F; // jal x0, 0
        */
        /*
        // 1. LUI (Load Upper Immediate)
        // [PC=0] rom[0]: lui x10, 0xABCDE
        // 예상 결과: x10 = 0xABCDE000 (imm을 12비트 왼쪽 시프트)
        rom[0] = 32'hABCDE537;

        // 2. AUIPC (Add Upper Immediate to PC)
        // [PC=4] rom[1]: auipc x11, 0x12345
        // 예상 결과: x11 = PC + (0x12345 << 12) = 4 + 0x12345000 = 0x12345004
        rom[1] = 32'h12345597;

        // 3. JAL (Jump and Link)
        // [PC=8] rom[2]: jal x12, 8 (PC + 8 = 16, 즉 rom[4]로 점프)
        // 예상 결과: x12 = PC + 4 = 12 (복귀 주소 저장)
        // PC는 rom[3]을 건너뛰고 16 (rom[4]의 주소)이 됨
        rom[2] = 32'h0080066F; // J-Type encoding for imm=8

        // 4. SKIPPED
        // [PC=12] rom[3]: (rom[2]의 JAL에 의해 실행되지 않음)
        rom[3] = 32'hDEADBEEF; // JAL이 실패하면 이 명령어가 실행됨

        // 5. JALR (Jump and Link Register)
        // [PC=16] rom[4]: jalr x13, x1, 19 (rs1=x1=1, imm=19)
        // 점프 타겟: (x1 + 19) = 1 + 19 = 20 (rom[5]의 주소)
        // 예상 결과: x13 = PC + 4 = 16 + 4 = 20 (복귀 주소 저장)
        // PC는 20 (rom[5]의 주소)이 됨
        rom[4] = 32'h013086E7; // I-Type encoding for JALR

        // 6. 테스트 종료 (무한 루프)
        // [PC=20] rom[5]: jal x0, 0 (현재 위치로 점프)
        rom[5] = 32'h0000006F;
         */
         /*
        // --- 1. 테스트 값 설정 ---
        // x5 = -100 (0xFFFFFF9C)
        rom[0] = 32'hF9C00293; // addi x5, x0, -100

        // --- 2. S-Type (Store) : x0(0번지) 기준으로 저장 ---
        // Mem[4] = 0xFFFFFF9C (Word)
        rom[1] = 32'h00502223; // sw x5, 4(x0)
        
        // Mem[8] = 0xFF9C (Half-word)
        rom[2] = 32'h00501423; // sh x5, 8(x0)
        
        // Mem[12] = 0x9C (Byte)
        rom[3] = 32'h00500623; // sb x5, 12(x0)

        // --- 3. L-Type (Load) : x0(0번지) 기준으로 로드 ---
        // LW: x10 = Mem[4]
        rom[4] = 32'h00402503; // lw x10, 4(x0)
        
        // LH: x11 = Mem[8] (부호 확장)
        rom[5] = 32'h00801583; // lh x11, 8(x0)
        
        // LHU: x12 = Mem[8] (0으로 확장)
        rom[6] = 32'h00805603; // lhu x12, 8(x0)
        
        // LB: x13 = Mem[12] (부호 확장)
        rom[7] = 32'h00C00683; // lb x13, 12(x0)
        
        // LBU: x14 = Mem[12] (0으로 확장)
        rom[8] = 32'h00C04703; // lbu x14, 12(x0)

        // --- 4. 테스트 종료 ---
        rom[9] = 32'h0000006F; // jal x0, 0 (무한 루프)
        */

        // //rom[x]=32'b   f7  _ rs2 _ rs1 _ f3_ rd  _ opcode;// R-Type
        // rom[0] = 32'b0000000_00001_00010_000_00100_0110011;// add x4, x2, x1
        // rom[1] = 32'b0100000_00001_00010_000_00101_0110011;// sub x5, x2, x1
        // rom[2] = 32'b0000000_00000_00011_111_00110_0110011;// and x6, x3, x0
        // rom[3] = 32'b0000000_00000_00011_110_00111_0110011;// or  x7, x3, x0
        // //rom[x]=32'b   imm      _ rs1 _ f3_ rd  _ opcode; // I-Type
        // rom[4] = 32'b000000000001_00001_000_01001_0010011;// addi x9, x1, 1;
        // rom[5] = 32'b000000000100_00010_111_01010_0010011;// andi x10, x2, 4;
        // rom[6] = 32'b000000000011_00001_001_01011_0010011;// slli x11, x1, 3;
        // rom[7] = 32'b000000001001_00001_001_01100_0010011;// slli x12, x1, 9;
        // rom[8] = 32'b000000011110_00001_001_01101_0010011;// slli x13, x1, 30;
        // //rom[x]=32'b imm(7)_ rs2 _ rs1 _ f3_imm5 _ opcode; // B-Type
        // rom[9] = 32'b0000000_00010_00001_000_01000_1100011;// beq x1, x2, 8;
        // //rom[x]=32'b imm(7)_ rs2 _ rs1 _ f3_imm5 _ opcode; // S-Type
        // rom[10] = 32'b0000000_01011_00000_000_00100_0100011;// sb x11, 4(x0);
        // rom[11]= 32'b0000000_01100_00000_001_01000_0100011;// sh x12, 8(x0);
        // rom[12]= 32'b0000000_01101_00000_010_01100_0100011;// sw x13, 12(x0);
        // //rom[x]=32'b    imm(12)  _ rs1 _ f3_ rd  _ opcode; // L-Type
        // rom[13] = 32'b000000000100_00000_000_01110_0000011;// lb x14, 4(x0);
        // rom[14] = 32'b000000001000_00000_001_01111_0000011;// lh x15, 8(x0);
        // rom[15] = 32'b000000001100_00000_010_10000_0000011;// lw x16, 12(x0);
        // //rom[x]=32'b    imm(20)            _ rd  _ opcode;// L-Type
        // rom[16] =   32'b00010000000000000000_10001_0110111;// lui x17, 0x10000000;
        
    end

    assign data = rom[addr[31:2]];
endmodule
